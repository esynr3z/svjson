class json_number extends json_value;
endclass : json_number