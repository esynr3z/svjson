class json_null extends json_value;
endclass : json_null