class json_string extends json_value;
endclass : json_string