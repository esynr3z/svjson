// Base JSON value
virtual class json_value;
    //pure virtual function json_value_e kind();
endclass : json_value
