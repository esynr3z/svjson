class json_array extends json_value;
endclass : json_array