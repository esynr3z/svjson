// Base JSON value
virtual class json_value;
endclass : json_value
