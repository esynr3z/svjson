// Generic interface for a class that can be encoded as JSON value
interface class json_value_encodable;
endclass : json_value_encodable
