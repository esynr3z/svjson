package json_pkg;

  // Forward declarations
  typedef json_value;
  typedef json_object;
  typedef json_array;
  typedef json_string;
  typedef json_int;
  typedef json_real;
  typedef json_bool;

  // Additional aliases for aggregate types
  typedef json_value json_value_queue_t[$];
  typedef json_value json_value_map_t[string];

  // All kinds of JSON value
  typedef enum {
    JSON_VALUE_OBJECT,
    JSON_VALUE_ARRAY,
    JSON_VALUE_STRING,
    JSON_VALUE_INT,
    JSON_VALUE_REAL,
    JSON_VALUE_BOOL
  } json_value_e;

  // Alias to raise syntax errors in a more compact way
  `define JSON_SYNTAX_ERR(KIND, STR, IDX, DESCR="")\
    parser_result::err( \
      json_error::create( \
        .kind(KIND), \
        .description(DESCR), \
        .json_str(STR), \
        .json_idx(IDX), \
        .source_file(`__FILE__), \
        .source_line(`__LINE__) \
      ) \
    )

  // Alias to raise internal error in a more compact way
  `define JSON_INTERNAL_ERR(DESCR="")\
    parser_result::err( \
      json_error::create( \
        .kind(json_error::INTERNAL), \
        .description(DESCR), \
        .source_file(`__FILE__), \
        .source_line(`__LINE__) \
      ) \
    )

  `include "json_error.sv"
  `include "json_result.sv"
  `include "json_value.sv"
  `include "json_object.sv"
  `include "json_array.sv"
  `include "json_string.sv"
  `include "json_int.sv"
  `include "json_real.sv"
  `include "json_bool.sv"

  `include "json_decoder.sv"

  `undef JSON_SYNTAX_ERR
  `undef JSON_INTERNAL_ERR
endpackage : json_pkg
