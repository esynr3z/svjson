class json_bool extends json_value;
endclass : json_bool