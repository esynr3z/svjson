class json_object extends json_value;
  json_value values[string];
endclass : json_object
