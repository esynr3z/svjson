package json_pkg;

endpackage : json_pkg
