package test_utils_pkg;
endpackage : test_utils_pkg